

module tb;

  reg clk;

  initial clk = 1'b1;

  always #10 clk = !clk;


  reg a, b, clear;

  wire r

  serial_adder #(.W(8)) adder(

  );

endmodule
