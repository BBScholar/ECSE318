

module mux8x1 #(parameter W = 8) (
  input [W-1:0] a, b, c, d, e, f, g, h,
  input sel,
  output [W-1:0] z
);




endmodule
