


module sign_extend
#(
  parameter IW=8,
  parameter OW=8
)
();


endmodule
